LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_arith.ALL;
USE ieee.std_logic_unsigned.ALL;
USE std.textio.ALL;

ENTITY ImageTestbench IS PORT 
(
	 pixelclock_input		: IN  std_logic;
	 resetclock_input		: IN  std_logic;
	 framesync_input		: IN  std_logic;
	 rowsync_input		   : IN  std_logic;
	 pixeldata_input		: IN  std_logic_vector(7 DOWNTO 0);
	 columnsrgb_output	: OUT std_logic_vector(15 DOWNTO 0);
	 rowsrgb_output		: OUT std_logic_vector(15 DOWNTO 0);
	 columnsgray_output	: OUT std_logic_vector(15 DOWNTO 0);
	 rowsgray_output		: OUT std_logic_vector(15 DOWNTO 0);
	 rowsync_output		: OUT std_logic;
	 framesync_output		: OUT std_logic;
	 pixeldata_output		: OUT std_logic_vector(7 DOWNTO 0) 
);		 
END ImageTestbench;

ARCHITECTURE behavioral OF ImageTestbench IS	
 
	TYPE ByteT IS (c0,c1,c2,c3,c4,c5,c6,c7,c8,c9,c10,c11,c12,c13,c14,c15,c16,c17,c18,
						c19,c20,c21,c22,c23,c24,c25,c26,c27,c28,c29,c30,c31,c32,c33,c34,
						c35,c36,c37,c38,c39,c40,c41,c42,c43,c44,c45,c46,c47,c48,c49,c50,
						c51,c52,c53,c54,c55,c56,c57,c58,c59,c60,c61,c62,c63,c64,c65,c66,
						c67,c68,c69,c70,c71,c72,c73,c74,c75,c76,c77,c78,c79,c80,c81,c82,
						c83,c84,c85,c86,c87,c88,c89,c90,c91,c92,c93,c94,c95,c96,c97,c98,
						c99,c100,c101,c102,c103,c104,c105,c106,c107,c108,c109,c110,c111,
						c112,c113,c114,c115,c116,c117,c118,c119,c120,c121,c122,c123,c124,
						c125,c126,c127,c128,c129,c130,c131,c132,c133,c134,c135,c136,c137,
						c138,c139,c140,c141,c142,c143,c144,c145,c146,c147,c148,c149,c150,
						c151,c152,c153,c154,c155,c156,c157,c158,c159,c160,c161,c162,c163,
						c164,c165,c166,c167,c168,c169,c170,c171,c172,c173,c174,c175,c176,
						c177,c178,c179,c180,c181,c182,c183,c184,c185,c186,c187,c188,c189,
						c190,c191,c192,c193,c194,c195,c196,c197,c198,c199,c200,c201,c202,
						c203,c204,c205,c206,c207,c208,c209,c210,c211,c212,c213,c214,c215,
						c216,c217,c218,c219,c220,c221,c222,c223,c224,c225,c226,c227,c228,
						c229,c230,c231,c232,c233,c234,c235,c236,c237,c238,c239,c240,c241,
				c242,c243,c244,c245,c246,c247,c248,c249,c250,c251,c252,c253,c254,c255);
  SUBTYPE Byte IS ByteT;
  TYPE ByteFileType IS FILE OF Byte;
  FILE infile	: ByteFileType OPEN read_mode IS "test1.bmp";
  FILE outfile	: ByteFileType OPEN write_mode IS "result.bmp";
    
  -- integer to bit_vector conversion
  
  FUNCTION int2bit_vec(A: integer; SIZE: integer) RETURN bit_vector IS
	VARIABLE RESULT: bit_vector(SIZE-1 DOWNTO 0);
	VARIABLE TMP	: integer;
	BEGIN
		TMP := A;
		FOR i IN 0 TO SIZE - 1 LOOP
			IF TMP mod 2 = 1 THEN RESULT(i) := '1';
			ELSE RESULT(i) := '0';
			END IF;
			TMP := TMP / 2;
		END LOOP;
		RETURN RESULT;
	END;

  BEGIN  

	read_image : PROCESS (pixelclock_input)
	VARIABLE pixelB 		: Byte;
	VARIABLE pixelG 		: Byte;
	VARIABLE pixelR 		: Byte;
	VARIABLE pixel_color : Byte;
	VARIABLE pixel_gray  : integer;
	VARIABLE columnsrgb	: std_logic_vector(15 DOWNTO 0);
	VARIABLE rowsrgb		: std_logic_vector(15 DOWNTO 0);
	VARIABLE columnsgray	: std_logic_vector(15 DOWNTO 0);
	VARIABLE rowsgray		: std_logic_vector(15 DOWNTO 0);
	VARIABLE count			: integer;
	VARIABLE rowsync		: std_logic := '0';
	VARIABLE framesync	: std_logic := '0';
	VARIABLE stop			: std_logic;
  
	BEGIN  -- PROCESS read_image
		IF (resetclock_input = '1') THEN
			pixeldata_output <= (OTHERS => '0');
			rowsync_output   <= '0';
			framesync_output <= '0';
			columnsgray	     := (OTHERS => '0');
			rowsgray		     := (OTHERS => '0');
		FOR i IN 0 to 53 LOOP -- read header infos
			read(infile, pixel_color);
			write(outfile, pixel_color);
			CASE i IS
				WHEN 18 => columnsrgb(7 DOWNTO 0)  := to_stdlogicvector(int2bit_vec(ByteT'POS(pixel_color), 8)); -- 1st byte of columnsrgb 
				WHEN 19 => columnsrgb(15 DOWNTO 8) := to_stdlogicvector(int2bit_vec(ByteT'POS(pixel_color), 8)); -- 2nd byte of columnsrgb
				WHEN 22 => rowsrgb(7 DOWNTO 0) 	  := to_stdlogicvector(int2bit_vec(ByteT'POS(pixel_color), 8)); -- 1st byte of rowsrgb
				WHEN 23 => rowsrgb(15 DOWNTO 8)    := to_stdlogicvector(int2bit_vec(ByteT'POS(pixel_color), 8)); -- 2nd byte of rowsrgb
				WHEN 24 => columnsrgb_output <= columnsrgb; rowsrgb_output	<= rowsrgb; columnsrgb := columnsrgb - 1; rowsrgb := rowsrgb - 1;
				WHEN OTHERS => NULL;
			END CASE;
		END LOOP; -- i
		rowsync   := '1';
		framesync := '1';
		count	    := 10;
		stop	    := '0';
		
		ELSIF (pixelclock_input'EVENT and pixelclock_input = '1') THEN	
		
			rowsync_output   <= rowsync;
			framesync_output <= framesync;
			
			IF rowsync = '1' THEN	
			
				IF stop = '0' THEN
					read(infile, pixelB); 
					read(infile, pixelG);
					read(infile, pixelR); 
					pixel_gray := (ByteT'POS(pixelB)*11) + (ByteT'POS(pixelR)*30) + (ByteT'POS(pixelG)*59);
					pixel_gray := pixel_gray / 100;
					pixeldata_output	 <= CONV_STD_LOGIC_VECTOR(integer(pixel_gray), 8);
					columnsgray_output <= columnsgray;
					rowsgray_output	 <= rowsgray;
					
				END IF;
				
				IF columnsgray = columnsrgb THEN
					columnsgray	:= (OTHERS => '0');
					rowsync	   := '0';
					IF rowsgray = rowsrgb THEN
						File_Close(infile);
						rowsgray	 := (OTHERS => '0');
						framesync := '0';
						stop      := '1';
					ELSE
						rowsgray := rowsgray + 1;
					END IF;		-- rowsgray
				ELSE
					columnsgray := columnsgray + 1;
				END IF;			-- columnsgray
				
			ELSE					-- rowsync
				IF count > 0 THEN
					count	:= count -1;
				ELSE
					count	    := 10;
					rowsync   := '1';
					framesync := '1';
				END IF;
				pixeldata_output <= (OTHERS => 'X');
			END IF;	-- rowsync
		
		IF framesync_input = '1' THEN
			IF rowsync_input = '1' THEN
				write(outfile, ByteT'VAL(ieee.numeric_std.to_Integer(ieee.numeric_std.unsigned(pixeldata_input)))); 				
				write(outfile, ByteT'VAL(ieee.numeric_std.to_Integer(ieee.numeric_std.unsigned(pixeldata_input)))); 
				write(outfile, ByteT'VAL(ieee.numeric_std.to_Integer(ieee.numeric_std.unsigned(pixeldata_input)))); 
			END IF; -- rowsync_input
		END IF; --frsync_i
	 END IF; -- clk
  END PROCESS read_image;
  
END behavioral;